module SBoxInv(in, out);
input wire[0:127]in;
output wire[0:127]out;
genvar i;
generate
for (i = 0; i < 127; i = i + 8)
	begin:hi
	assign out[i:i + 7] =
	(in[i:i+7] == 8'b 0110_0011) ? 8'b00000000:
(in[i:i+7] == 8'b 0111_1100) ? 8'b00000001:
(in[i:i+7] == 8'b 0111_0111) ? 8'b00000010:
(in[i:i+7] == 8'b 0111_1011) ? 8'b00000011 :
(in[i:i+7] == 8'b 1111_0010) ? 8'b00000100:
(in[i:i+7] == 8'b 0110_1011) ? 8'b00000101:
(in[i:i+7] == 8'b 0110_1111) ? 8'b00000110:
(in[i:i+7] == 8'b 1100_0101) ? 8'b00000111:
(in[i:i+7] == 8'b 0011_0000) ? 8'b00001000:
(in[i:i+7] == 8'b 0000_0001) ? 8'b00001001:
(in[i:i+7] == 8'b 0110_0111) ? 8'b00001010:
(in[i:i+7] == 8'b 0010_1011) ? 8'b00001011:
(in[i:i+7] == 8'b 1111_1110) ? 8'b00001100:
(in[i:i+7] == 8'b 1101_0111) ? 8'b00001101:
(in[i:i+7] == 8'b 1010_1011) ? 8'b00001110:
(in[i:i+7] == 8'b 0111_0110) ? 8'b00001111:

(in[i:i+7] == 8'b 1100_1010) ? 8'b00010000:
(in[i:i+7] == 8'b 1000_0010) ? 8'b00010001:
(in[i:i+7] == 8'b 1100_1001) ? 8'b00010010:
(in[i:i+7] == 8'b 0111_1101) ? 8'b00010011:
(in[i:i+7] == 8'b 1111_1010) ? 8'b00010100:
(in[i:i+7] == 8'b 0101_1001) ? 8'b00010101:
(in[i:i+7] == 8'b 0100_0111) ? 8'b00010110:
(in[i:i+7] == 8'b 1111_0000) ? 8'b00010111:
(in[i:i+7] == 8'b 1010_1101) ? 8'b00011000:
(in[i:i+7] == 8'b 1101_0100) ? 8'b00011001:
(in[i:i+7] == 8'b 1010_0010) ? 8'b00011010:
(in[i:i+7] == 8'b 1010_1111) ? 8'b00011011:
(in[i:i+7] == 8'b 1001_1100) ? 8'b00011100:
(in[i:i+7] == 8'b 1010_0100) ? 8'b00011101:
(in[i:i+7] == 8'b 0111_0010) ? 8'b00011110 :
(in[i:i+7] == 8'b 1100_0000) ? 8'b00011111:

(in[i:i+7] == 8'b 1011_0111) ? 8'b00100000:
(in[i:i+7] == 8'b 1111_1101) ? 8'b00100001:
(in[i:i+7] == 8'b 1001_0011) ? 8'b00100010:
(in[i:i+7] == 8'b 0010_0110) ? 8'b00100011:
(in[i:i+7] == 8'b 0011_0110) ? 8'b00100100:
(in[i:i+7] == 8'b 0011_1111) ? 8'b00100101:
(in[i:i+7] == 8'b 1111_0111) ? 8'b00100110:
(in[i:i+7] == 8'b 1100_1100) ? 8'b00100111:
(in[i:i+7] == 8'b 0011_0100) ? 8'b00101000:
(in[i:i+7] == 8'b 1010_0101) ? 8'b00101001:
(in[i:i+7] == 8'b 1110_0101) ? 8'b00101010:
(in[i:i+7] == 8'b 1111_0001) ? 8'b00101011:
(in[i:i+7] == 8'b 0111_0001) ? 8'b00101100:
(in[i:i+7] == 8'b 1101_1000) ? 8'b00101101:
(in[i:i+7] == 8'b 0011_0001) ? 8'b00101110:
(in[i:i+7] == 8'b 0001_0101) ? 8'b00101111:

(in[i:i+7] == 8'b 0000_0100) ? 8'b00110000:
(in[i:i+7] == 8'b 1100_0111) ? 8'b00110001:
(in[i:i+7] == 8'b 0010_0011) ? 8'b00110010:
(in[i:i+7] == 8'b 1100_0011) ? 8'b00110011:
(in[i:i+7] == 8'b 0001_1000) ? 8'b00110100:
(in[i:i+7] == 8'b 1001_0110) ? 8'b00110101:
(in[i:i+7] == 8'b 0000_0101) ? 8'b00110110:
(in[i:i+7] == 8'b 1001_1010) ? 8'b00110111:
(in[i:i+7] == 8'b 0000_0111) ? 8'b00111000:
(in[i:i+7] == 8'b 0001_0010) ? 8'b00111001:
(in[i:i+7] == 8'b 1000_0000) ? 8'b00111010:
(in[i:i+7] == 8'b 1110_0010) ? 8'b00111011:
(in[i:i+7] == 8'b 1110_1011) ? 8'b00111100:
(in[i:i+7] == 8'b 0010_0111) ? 8'b00111101:
(in[i:i+7] == 8'b 1011_0010) ? 8'b00111110:
(in[i:i+7] == 8'b 0111_0101) ? 8'b00111111:

(in[i:i+7] == 8'b 0000_1001) ? 8'b01000000:
(in[i:i+7] == 8'b 1000_0011) ? 8'b01000001:
(in[i:i+7] == 8'b 0010_1100) ? 8'b01000010:
(in[i:i+7] == 8'b 0001_1010) ? 8'b01000011:
(in[i:i+7] == 8'b 0001_1011) ? 8'b01000100:
(in[i:i+7] == 8'b 0110_1110) ? 8'b01000101:
(in[i:i+7] == 8'b 0101_1010) ? 8'b01000110:
(in[i:i+7] == 8'b 1010_0000) ? 8'b01000111:
(in[i:i+7] == 8'b 0101_0010) ? 8'b01001000:
(in[i:i+7] == 8'b 0011_1011) ? 8'b01001001:
(in[i:i+7] == 8'b 1101_0110) ? 8'b01001010:
(in[i:i+7] == 8'b 1011_0011) ? 8'b01001011:
(in[i:i+7] == 8'b 0010_1001) ? 8'b01001100:
(in[i:i+7] == 8'b 1110_0011) ? 8'b01001101:
(in[i:i+7] == 8'b 0010_1111) ? 8'b01001110:
(in[i:i+7] == 8'b 1000_0100) ? 8'b01001111:

(in[i:i+7] == 8'b 0101_0011) ? 8'b01010000:
(in[i:i+7] == 8'b 1101_0001) ? 8'b01010001:
(in[i:i+7] == 8'b 0000_0000) ? 8'b01010010:
(in[i:i+7] == 8'b 1110_1101) ? 8'b01010011:
(in[i:i+7] == 8'b 0010_0000) ? 8'b01010100:
(in[i:i+7] == 8'b 1111_1100) ? 8'b01010101:
(in[i:i+7] == 8'b 1011_0001) ? 8'b01010110:
(in[i:i+7] == 8'b 0101_1011) ? 8'b01010111:
(in[i:i+7] == 8'b 0110_1010) ? 8'b01011000:
(in[i:i+7] == 8'b 1100_1011) ? 8'b01011001:
(in[i:i+7] == 8'b 1011_1110) ? 8'b01011010:
(in[i:i+7] == 8'b 0011_1001) ? 8'b01011011:
(in[i:i+7] == 8'b 0100_1010) ? 8'b01011100:
(in[i:i+7] == 8'b 0100_1100) ? 8'b01011101:
(in[i:i+7] == 8'b 0101_1000) ? 8'b01011110:
(in[i:i+7] == 8'b 1100_1111) ? 8'b01011111:

(in[i:i+7] == 8'b 1101_0000) ? 8'b01100000:
(in[i:i+7] == 8'b 1110_1111) ? 8'b01100001:
(in[i:i+7] == 8'b 1010_1010) ? 8'b01100010:
(in[i:i+7] == 8'b 1111_1011) ? 8'b01100011:
(in[i:i+7] == 8'b 0100_0011) ? 8'b01100100:
(in[i:i+7] == 8'b 0100_1101) ? 8'b01100101:
(in[i:i+7] == 8'b 0011_0011) ? 8'b01100110:
(in[i:i+7] == 8'b 1000_0101) ? 8'b01100111:
(in[i:i+7] == 8'b 0100_0101) ? 8'b01101000:
(in[i:i+7] == 8'b 1111_1001) ? 8'b01101001:
(in[i:i+7] == 8'b 0000_0010) ? 8'b01101010:
(in[i:i+7] == 8'b 0111_1111) ? 8'b01101011:
(in[i:i+7] == 8'b 0101_0000) ? 8'b01101100:
(in[i:i+7] == 8'b 0011_1100) ? 8'b01101101:
(in[i:i+7] == 8'b 1001_1111) ? 8'b01101110:
(in[i:i+7] == 8'b 1010_1000) ? 8'b01101111:

(in[i:i+7] == 8'b 0101_0001) ? 8'b01110000:
(in[i:i+7] == 8'b 1010_0011) ? 8'b01110001:
(in[i:i+7] == 8'b 0100_0000) ? 8'b01110010:
(in[i:i+7] == 8'b 1000_1111) ? 8'b01110011:
(in[i:i+7] == 8'b 1001_0010) ? 8'b01110100:
(in[i:i+7] == 8'b 1001_1101) ? 8'b01110101:
(in[i:i+7] == 8'b 0011_1000) ? 8'b01110110:
(in[i:i+7] == 8'b 1111_0101) ? 8'b01110111:
(in[i:i+7] == 8'b 1011_1100) ? 8'b01111000:
(in[i:i+7] == 8'b 1011_0110) ? 8'b01111001:
(in[i:i+7] == 8'b 1101_1010) ? 8'b01111010:
(in[i:i+7] == 8'b 0010_0001) ? 8'b01111011:
(in[i:i+7] == 8'b 0001_0000) ? 8'b01111100:
(in[i:i+7] == 8'b 1111_1111) ? 8'b01111101:
(in[i:i+7] == 8'b 1111_0011) ? 8'b01111110:
(in[i:i+7] == 8'b 1101_0010) ? 8'b01111111:

(in[i:i+7] == 8'b 1100_1101) ? 8'b10000000:
(in[i:i+7] == 8'b 0000_1100) ? 8'b10000001:
(in[i:i+7] == 8'b 0001_0011) ? 8'b10000010:
(in[i:i+7] == 8'b 1110_1100) ? 8'b10000011:
(in[i:i+7] == 8'b 0101_1111) ? 8'b10000100:
(in[i:i+7] == 8'b 1001_0111) ? 8'b10000101:
(in[i:i+7] == 8'b 0100_0100) ? 8'b10000110:
(in[i:i+7] == 8'b 0001_0111) ? 8'b10000111:
(in[i:i+7] == 8'b 1100_0100) ? 8'b10001000:
(in[i:i+7] == 8'b 1010_0111) ? 8'b10001001:
(in[i:i+7] == 8'b 0111_1110) ? 8'b10001010:
(in[i:i+7] == 8'b 0011_1101) ? 8'b10001011:
(in[i:i+7] == 8'b 0110_0100) ? 8'b10001100:
(in[i:i+7] == 8'b 0101_1101) ? 8'b10001101:
(in[i:i+7] == 8'b 0001_1001) ? 8'b10001110:
(in[i:i+7] == 8'b 0111_0011) ? 8'b10001111:

(in[i:i+7] == 8'b 0110_0000) ? 8'b10010000:
(in[i:i+7] == 8'b 1000_0001) ? 8'b10010001:
(in[i:i+7] == 8'b 0100_1111) ? 8'b10010010:
(in[i:i+7] == 8'b 1101_1100) ? 8'b10010011:
(in[i:i+7] == 8'b 0010_0010) ? 8'b10010100:
(in[i:i+7] == 8'b 0010_1010) ? 8'b10010101:
(in[i:i+7] == 8'b 1001_0000) ? 8'b10010110:
(in[i:i+7] == 8'b 1000_1000) ? 8'b10010111:
(in[i:i+7] == 8'b 0100_0110) ? 8'b10011000:
(in[i:i+7] == 8'b 1110_1110) ? 8'b10011001:
(in[i:i+7] == 8'b 1011_1000) ? 8'b10011010:
(in[i:i+7] == 8'b 0001_0100) ? 8'b10011011:
(in[i:i+7] == 8'b 1101_1110) ? 8'b10011100:
(in[i:i+7] == 8'b 0101_1110) ? 8'b10011101:
(in[i:i+7] == 8'b 0000_1011) ? 8'b10011110:
(in[i:i+7] == 8'b 1101_1011) ? 8'b10011111:

(in[i:i+7] == 8'b 1110_0000) ? 8'b10100000:
(in[i:i+7] == 8'b 0011_0010) ? 8'b10100001:
(in[i:i+7] == 8'b 0011_1010) ? 8'b10100010:
(in[i:i+7] == 8'b 0000_1010) ? 8'b10100011:
(in[i:i+7] == 8'b 0100_1001) ? 8'b10100100:
(in[i:i+7] == 8'b 0000_0110) ? 8'b10100101:
(in[i:i+7] == 8'b 0010_0100) ? 8'b10100110:
(in[i:i+7] == 8'b 0101_1100) ? 8'b10100111:
(in[i:i+7] == 8'b 1100_0010) ? 8'b10101000:
(in[i:i+7] == 8'b 1101_0011) ? 8'b10101001:
(in[i:i+7] == 8'b 1010_1100) ? 8'b10101010:
(in[i:i+7] == 8'b 0110_0010) ? 8'b10101011:
(in[i:i+7] == 8'b 1001_0001) ? 8'b10101100:
(in[i:i+7] == 8'b 1001_0101) ? 8'b10101101:
(in[i:i+7] == 8'b 1110_0100) ? 8'b10101110:
(in[i:i+7] == 8'b 0111_1001) ? 8'b10101111:

(in[i:i+7] == 8'b 1110_0111) ? 8'b10110000:
(in[i:i+7] == 8'b 1100_1000) ? 8'b10110001:
(in[i:i+7] == 8'b 0011_0111) ? 8'b10110010:
(in[i:i+7] == 8'b 0110_1101) ? 8'b10110011:
(in[i:i+7] == 8'b 1000_1101) ? 8'b10110100:
(in[i:i+7] == 8'b 1101_0101) ? 8'b10110101:
(in[i:i+7] == 8'b 0100_1110) ? 8'b10110110:
(in[i:i+7] == 8'b 1010_1001) ? 8'b10110111:
(in[i:i+7] == 8'b 0110_1100) ? 8'b10111000:
(in[i:i+7] == 8'b 0101_0110) ? 8'b10111001:
(in[i:i+7] == 8'b 1111_0100) ? 8'b10111010:
(in[i:i+7] == 8'b 1110_1010) ? 8'b10111011:
(in[i:i+7] == 8'b 0110_0101) ? 8'b10111100:
(in[i:i+7] == 8'b 0111_1010) ? 8'b10111101:
(in[i:i+7] == 8'b 1010_1110) ? 8'b10111110:
(in[i:i+7] == 8'b 0000_1000) ? 8'b10111111:

(in[i:i+7] == 8'b 1011_1010) ? 8'b11000000:
(in[i:i+7] == 8'b 0111_1000) ? 8'b11000001:
(in[i:i+7] == 8'b 0010_0101) ? 8'b11000010:
(in[i:i+7] == 8'b 0010_1110) ? 8'b11000011:
(in[i:i+7] == 8'b 0001_1100) ? 8'b11000100:
(in[i:i+7] == 8'b 1010_0110) ? 8'b11000101:
(in[i:i+7] == 8'b 1011_0100) ? 8'b11000110:
(in[i:i+7] == 8'b 1100_0110) ? 8'b11000111:
(in[i:i+7] == 8'b 1110_1000) ? 8'b11001000:
(in[i:i+7] == 8'b 1101_1101) ? 8'b11001001:
(in[i:i+7] == 8'b 0111_0100) ? 8'b11001010:
(in[i:i+7] == 8'b 0001_1111) ? 8'b11001011:
(in[i:i+7] == 8'b 0100_1011) ? 8'b11001100:
(in[i:i+7] == 8'b 1011_1101) ? 8'b11001101:
(in[i:i+7] == 8'b 1000_1011) ? 8'b11001110:
(in[i:i+7] == 8'b 1000_1010) ? 8'b11001111:

(in[i:i+7] == 8'b 0111_0000) ? 8'b11010000:
(in[i:i+7] == 8'b 0011_1110) ? 8'b11010001:
(in[i:i+7] == 8'b 1011_0101) ? 8'b11010010:
(in[i:i+7] == 8'b 0110_0110) ? 8'b11010011:
(in[i:i+7] == 8'b 0100_1000) ? 8'b11010100:
(in[i:i+7] == 8'b 0000_0011) ? 8'b11010101:
(in[i:i+7] == 8'b 1111_0110) ? 8'b11010110:
(in[i:i+7] == 8'b 0000_1110) ? 8'b11010111:
(in[i:i+7] == 8'b 0110_0001) ? 8'b11011000:
(in[i:i+7] == 8'b 0011_0101) ? 8'b11011001:
(in[i:i+7] == 8'b 0101_0111) ? 8'b11011010:
(in[i:i+7] == 8'b 1011_1001) ? 8'b11011011:
(in[i:i+7] == 8'b 1000_0110) ? 8'b11011100:
(in[i:i+7] == 8'b 1100_0001) ? 8'b11011101:
(in[i:i+7] == 8'b 0001_1101) ? 8'b11011110:
(in[i:i+7] == 8'b 1001_1110) ? 8'b11011111:

(in[i:i+7] == 8'b 1110_0001) ? 8'b11100000:
(in[i:i+7] == 8'b 1111_1000) ? 8'b11100001:
(in[i:i+7] == 8'b 1001_1000) ? 8'b11100010:
(in[i:i+7] == 8'b 0001_0001) ? 8'b11100011:
(in[i:i+7] == 8'b 0110_1001) ? 8'b11100100:
(in[i:i+7] == 8'b 1101_1001) ? 8'b11100101:
(in[i:i+7] == 8'b 1000_1110) ? 8'b11100110:
(in[i:i+7] == 8'b 1001_0100) ? 8'b11100111:
(in[i:i+7] == 8'b 1001_1011) ? 8'b11101000:
(in[i:i+7] == 8'b 0001_1110) ? 8'b11101001:
(in[i:i+7] == 8'b 1000_0111) ? 8'b11101010:
(in[i:i+7] == 8'b 1110_1001) ? 8'b11101011:
(in[i:i+7] == 8'b 1100_1110) ? 8'b11101100:
(in[i:i+7] == 8'b 0101_0101) ? 8'b11101101:
(in[i:i+7] == 8'b 0010_1000) ? 8'b11101110:
(in[i:i+7] == 8'b 1101_1111) ? 8'b11101111:

(in[i:i+7] == 8'b 1000_1100) ? 8'b11110000:
(in[i:i+7] == 8'b 1010_0001) ? 8'b11110001:
(in[i:i+7] == 8'b 1000_1001) ? 8'b11110010:
(in[i:i+7] == 8'b 0000_1101) ? 8'b11110011:
(in[i:i+7] == 8'b 1011_1111) ? 8'b11110100:
(in[i:i+7] == 8'b 1110_0110) ? 8'b11110101:
(in[i:i+7] == 8'b 0100_0010) ? 8'b11110110:
(in[i:i+7] == 8'b 0110_1000) ? 8'b11110111:
(in[i:i+7] == 8'b 0100_0001) ? 8'b11111000:
(in[i:i+7] == 8'b 1001_1001) ? 8'b11111001:
(in[i:i+7] == 8'b 0010_1101) ? 8'b11111010:
(in[i:i+7] == 8'b 0000_1111) ? 8'b11111011:
(in[i:i+7] == 8'b 1011_0000) ? 8'b11111100:
(in[i:i+7] == 8'b 0101_0100) ? 8'b11111101:
(in[i:i+7] == 8'b 1011_1011) ? 8'b11111110:
(in[i:i+7] == 8'b 0001_0110) ? 8'b11111111:

8'bxxxxxxxx;
end
endgenerate
endmodule